`include "Slave.v"
module Master (

);


endmodule
