module Cipher #(parameter Nk = 4, parameter Nr = 10)(
                input [127:0] in,
                input [Nk*32 - 1:0] key,
                output [128 * (Nr + 1) - 1:0] key_out,
                output [127:0] out
);

wire [127:0] start [0:Nr];
wire [127:0] s_box [0:Nr - 1];
wire [127:0] s_row [0:Nr - 1];
wire [127:0] m_col [0:Nr - 1];
wire [127:0] k_sch [0:Nr];
wire [Nk*32*11 - 1:0] keys;
wire [128 * (Nr + 1) - 1:0] key_o;
wire [31:0] Rcon  [0:9];
assign Rcon[0] = 32'h01000000;
assign Rcon[1] = 32'h02000000;
assign Rcon[2] = 32'h04000000;
assign Rcon[3] = 32'h08000000;
assign Rcon[4] = 32'h10000000;
assign Rcon[5] = 32'h20000000;
assign Rcon[6] = 32'h40000000;
assign Rcon[7] = 32'h80000000;
assign Rcon[8] = 32'h1B000000;
assign Rcon[9] = 32'h36000000;


AddRoundKey add_key_strt (in, key[Nk*32 - 1 -: 128], start[0]);
assign keys[Nk*32*11 - 1 -: Nk*32] = key;

genvar i;
generate
    for (i = 0; i < 10; i = i + 1) begin : exp
        KeyExpansion #(Nk) key_exp (keys[Nk*32*(11 - i) - 1 -: Nk*32], Rcon[i][31:0], keys[Nk*32*(10 - i) - 1 -: Nk*32]);
    end
    for (i = 0; i <= Nr; i = i + 1) begin : to_block
        assign k_sch[i] = keys[Nk*32*11 - 1 - 128*i -: 128];
    end
    for (i = 0; i < Nr - 1; i = i + 1) begin : sim
        SubBytes sbox(start[i], s_box[i]);
        ShiftRows shift_rows(s_box[i], s_row[i]);
        MixColumns mix_col(s_row[i], m_col[i]);
        AddRoundKey add_key (m_col[i], k_sch[i + 1], start[i + 1]);
    end
endgenerate

SubBytes sbox(start[Nr - 1], s_box[Nr - 1]);
ShiftRows shift_rows(s_box[Nr - 1], s_row[Nr - 1]);
AddRoundKey add_key_end (s_row[Nr - 1], k_sch[Nr], start[Nr]);

generate
    for (i = 0; i <= Nr; i = i + 1) begin : to_line
       assign key_o [(128 *(Nr + 1 - i) - 1) -: 128] = k_sch[Nr - i];
    end
endgenerate

assign out = start[Nr];
assign key_out = key_o;

endmodule
